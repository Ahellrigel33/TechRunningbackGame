`timescale 1 ps / 1 ps
module rw_manager_m10_inst_ROM (
	clock,
	rdaddress,
	q);
	
	input	  clock;
	input	[6:0]  rdaddress;
	output	[19:0]  q;
	
	reg	[19:0]  q;
	
	wire	[6:0]  rdaddress_r;
  assign  rdaddress_r =   rdaddress;
	
always @ (posedge clock)
    case(rdaddress_r)
'h00 : q <= 'h080180;
'h01 : q <= 'h000100;
'h02 : q <= 'h080000;
'h03 : q <= 'h000200;
'h04 : q <= 'h080000;
'h05 : q <= 'h000280;
'h06 : q <= 'h080000;
'h07 : q <= 'h000300;
'h08 : q <= 'h080000;
'h09 : q <= 'h000380;
'h0A : q <= 'h080000;
'h0B : q <= 'h000400;
'h0C : q <= 'h080000;
'h0D : q <= 'h000480;
'h0E : q <= 'h080000;
'h0F : q <= 'h000500;
'h10 : q <= 'h080000;
'h11 : q <= 'h000600;
'h12 : q <= 'h008000;
'h13 : q <= 'h000680;
'h14 : q <= 'h00A000;
'h15 : q <= 'h080000;
'h16 : q <= 'h000700;
'h17 : q <= 'h080000;
'h18 : q <= 'h000780;
'h19 : q <= 'h080000;
'h1A : q <= 'h000968;
'h1B : q <= 'h00CAE8;
'h1C : q <= 'h0008E8;
'h1D : q <= 'h008AE8;
'h1E : q <= 'h000988;
'h1F : q <= 'h00EA88;
'h20 : q <= 'h000808;
'h21 : q <= 'h00AA88;
'h22 : q <= 'h080000;
'h23 : q <= 'h00CC00;
'h24 : q <= 'h00CB80;
'h25 : q <= 'h00E080;
'h26 : q <= 'h000A00;
'h27 : q <= 'h020AE0;
'h28 : q <= 'h020AE0;
'h29 : q <= 'h000B00;
'h2A : q <= 'h000000;
'h2B : q <= 'h000000;
'h2C : q <= 'h060C80;
'h2D : q <= 'h060E80;
'h2E : q <= 'h00A000;
'h2F : q <= 'h008000;
'h30 : q <= 'h080000;
'h31 : q <= 'h00CC00;
'h32 : q <= 'h00CB80;
'h33 : q <= 'h00E080;
'h34 : q <= 'h000A00;
'h35 : q <= 'h030AE0;
'h36 : q <= 'h030AE0;
'h37 : q <= 'h000B00;
'h38 : q <= 'h000000;
'h39 : q <= 'h000000;
'h3A : q <= 'h070C80;
'h3B : q <= 'h070E80;
'h3C : q <= 'h00A000;
'h3D : q <= 'h008000;
'h3E : q <= 'h080000;
'h3F : q <= 'h000F58;
'h40 : q <= 'h000058;
'h41 : q <= 'h080000;
'h42 : q <= 'h040C88;
'h43 : q <= 'h040E88;
'h44 : q <= 'h040D68;
'h45 : q <= 'h040EE8;
'h46 : q <= 'h00A000;
'h47 : q <= 'h040DE8;
'h48 : q <= 'h040EE8;
'h49 : q <= 'h040E08;
'h4A : q <= 'h040E88;
'h4B : q <= 'h000F00;
'h4C : q <= 'h00C000;
'h4D : q <= 'h008000;
'h4E : q <= 'h00E000;
'h4F : q <= 'h080000;
'h50 : q <= 'h000180;
'h51 : q <= 'h000180;
'h52 : q <= 'h00A180;
'h53 : q <= 'h008180;
'h54 : q <= 'h080180;
'h55 : q <= 'h008000;
'h56 : q <= 'h00A000;
'h57 : q <= 'h080000;
'h58 : q <= 'h000000;
'h59 : q <= 'h000000;
'h5A : q <= 'h000000;
'h5B : q <= 'h000000;
'h5C : q <= 'h000000;
'h5D : q <= 'h000000;
'h5E : q <= 'h000000;
'h5F : q <= 'h000000;
'h60 : q <= 'h000000;
'h61 : q <= 'h000000;
'h62 : q <= 'h000000;
'h63 : q <= 'h000000;
'h64 : q <= 'h000000;
'h65 : q <= 'h000000;
'h66 : q <= 'h000000;
'h67 : q <= 'h000000;
'h68 : q <= 'h000000;
'h69 : q <= 'h000000;
'h6A : q <= 'h000000;
'h6B : q <= 'h000000;
'h6C : q <= 'h000000;
'h6D : q <= 'h000000;
'h6E : q <= 'h000000;
'h6F : q <= 'h000000;
'h70 : q <= 'h000000;
'h71 : q <= 'h000000;
'h72 : q <= 'h000000;
'h73 : q <= 'h000000;
'h74 : q <= 'h000000;
'h75 : q <= 'h000000;
'h76 : q <= 'h000000;
'h77 : q <= 'h000000;
'h78 : q <= 'h000000;
'h79 : q <= 'h000000;
'h7A : q <= 'h000000;
'h7B : q <= 'h000000;
'h7C : q <= 'h000000;
'h7D : q <= 'h000000;
'h7E : q <= 'h000000;
'h7F : q <= 'h000000;
        default : q <= 0;
    endcase
endmodule
