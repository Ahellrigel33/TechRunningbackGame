-- SDRAM_ADR.VHD (a peripheral module for SCOMP)
-- 2020.10.25
--
-- This module controls the address selection of the SDRAM memory on the rising edge of CS.


LIBRARY IEEE;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE LPM.LPM_COMPONENTS.ALL;


ENTITY SDRAM_ADR IS
  PORT(
    RESETN      : IN  STD_LOGIC;
    CS          : IN  STD_LOGIC;
    ADDRESS_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    ADDRESS_IN  : IN  STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END SDRAM_ADR;


ARCHITECTURE a OF SDRAM_ADR IS
  BEGIN
    PROCESS (RESETN, CS)
      BEGIN
        IF (RESETN = '0') THEN
          ADDRESS_OUT <= x"0000";
        ELSIF (RISING_EDGE(CS)) THEN
          ADDRESS_OUT <= ADDRESS_IN;
        END IF;
      END PROCESS;
  END a;